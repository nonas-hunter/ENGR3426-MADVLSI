magic
tech sky130A
timestamp 1694404404
<< nwell >>
rect -140 -70 130 70
<< nmos >>
rect -20 -205 -5 -105
rect 20 -205 35 -105
<< pmos >>
rect -20 -50 -5 50
rect 45 -50 60 50
<< ndiff >>
rect -70 -120 -20 -105
rect -70 -190 -55 -120
rect -35 -190 -20 -120
rect -70 -205 -20 -190
rect -5 -205 20 -105
rect 35 -120 85 -105
rect 35 -190 50 -120
rect 70 -190 85 -120
rect 35 -205 85 -190
<< pdiff >>
rect -70 35 -20 50
rect -70 -35 -55 35
rect -35 -35 -20 35
rect -70 -50 -20 -35
rect -5 35 45 50
rect -5 -35 10 35
rect 30 -35 45 35
rect -5 -50 45 -35
rect 60 35 110 50
rect 60 -35 75 35
rect 95 -35 110 35
rect 60 -50 110 -35
<< ndiffc >>
rect -55 -190 -35 -120
rect 50 -190 70 -120
<< pdiffc >>
rect -55 -35 -35 35
rect 10 -35 30 35
rect 75 -35 95 35
<< psubdiff >>
rect -120 -120 -70 -105
rect -120 -190 -105 -120
rect -85 -190 -70 -120
rect -120 -205 -70 -190
<< nsubdiff >>
rect -120 35 -70 50
rect -120 -35 -105 35
rect -85 -35 -70 35
rect -120 -50 -70 -35
<< psubdiffcont >>
rect -105 -190 -85 -120
<< nsubdiffcont >>
rect -105 -35 -85 35
<< poly >>
rect -20 50 -5 65
rect 45 50 60 65
rect -20 -105 -5 -50
rect 45 -70 60 -50
rect 20 -85 60 -70
rect 20 -105 35 -85
rect -20 -220 -5 -205
rect -45 -230 -5 -220
rect -45 -250 -35 -230
rect -15 -250 -5 -230
rect -45 -260 -5 -250
rect 20 -220 35 -205
rect 20 -230 60 -220
rect 20 -250 30 -230
rect 50 -250 60 -230
rect 20 -260 60 -250
<< polycont >>
rect -35 -250 -15 -230
rect 30 -250 50 -230
<< locali >>
rect -115 35 -25 45
rect -115 -35 -105 35
rect -85 -35 -55 35
rect -35 -35 -25 35
rect -115 -45 -25 -35
rect 0 35 40 45
rect 0 -35 10 35
rect 30 -35 40 35
rect 0 -45 40 -35
rect 65 35 105 45
rect 65 -35 75 35
rect 95 -35 105 35
rect 65 -45 105 -35
rect 20 -110 40 -45
rect -115 -120 -25 -110
rect -115 -190 -105 -120
rect -85 -190 -55 -120
rect -35 -190 -25 -120
rect 20 -120 80 -110
rect 20 -130 50 -120
rect -115 -200 -25 -190
rect 40 -190 50 -130
rect 70 -180 80 -120
rect 70 -190 100 -180
rect 40 -200 100 -190
rect 80 -220 100 -200
rect -140 -230 -5 -220
rect -140 -240 -35 -230
rect -45 -250 -35 -240
rect -15 -250 -5 -230
rect -45 -260 -5 -250
rect 20 -230 60 -220
rect 20 -250 30 -230
rect 50 -250 60 -230
rect 80 -240 130 -220
rect 20 -260 60 -250
rect 20 -280 40 -260
rect -140 -300 40 -280
<< viali >>
rect -105 -35 -85 35
rect -55 -35 -35 35
rect 75 -35 95 35
rect -105 -190 -85 -120
rect -55 -190 -35 -120
<< metal1 >>
rect -140 35 130 45
rect -140 -35 -105 35
rect -85 -35 -55 35
rect -35 -35 75 35
rect 95 -35 130 35
rect -140 -45 130 -35
rect -140 -120 130 -110
rect -140 -190 -105 -120
rect -85 -190 -55 -120
rect -35 -190 130 -120
rect -140 -200 130 -190
<< labels >>
rlabel locali -140 -230 -140 -230 7 A
port 1 w
rlabel locali -140 -290 -140 -290 7 B
port 2 w
rlabel locali 130 -230 130 -230 3 Y
port 3 e
rlabel metal1 -140 0 -140 0 7 VP
port 4 w
rlabel metal1 -140 -155 -140 -155 7 VN
port 5 w
<< end >>
