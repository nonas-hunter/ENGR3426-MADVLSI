magic
tech sky130A
timestamp 1695979802
<< nwell >>
rect -85 430 250 945
<< nmos >>
rect -20 -15 -5 385
rect 35 285 50 385
rect 100 285 115 385
rect 165 285 180 385
rect 35 -15 50 85
rect 100 -15 115 85
rect 165 -15 180 85
<< pmos >>
rect -20 745 -5 845
rect 50 745 65 845
rect -20 450 -5 550
rect 50 450 65 550
rect 115 450 130 845
rect 165 745 180 845
rect 165 450 180 550
<< ndiff >>
rect -65 370 -20 385
rect -65 300 -55 370
rect -35 300 -20 370
rect -65 285 -20 300
rect -45 85 -20 285
rect -65 70 -20 85
rect -65 0 -55 70
rect -35 0 -20 70
rect -65 -15 -20 0
rect -5 285 35 385
rect 50 370 100 385
rect 50 300 65 370
rect 85 300 100 370
rect 50 285 100 300
rect 115 370 165 385
rect 115 300 130 370
rect 150 300 165 370
rect 115 285 165 300
rect 180 370 230 385
rect 180 300 195 370
rect 215 300 230 370
rect 180 285 230 300
rect -5 85 25 285
rect -5 -15 35 85
rect 50 70 100 85
rect 50 0 65 70
rect 85 0 100 70
rect 50 -15 100 0
rect 115 70 165 85
rect 115 0 130 70
rect 150 0 165 70
rect 115 -15 165 0
rect 180 70 230 85
rect 180 0 195 70
rect 215 0 230 70
rect 180 -15 230 0
<< pdiff >>
rect -65 830 -20 845
rect -65 760 -55 830
rect -35 760 -20 830
rect -65 745 -20 760
rect -5 830 50 845
rect -5 760 10 830
rect 35 760 50 830
rect -5 745 50 760
rect 65 830 115 845
rect 65 760 80 830
rect 100 760 115 830
rect 65 745 115 760
rect 90 550 115 745
rect -65 535 -20 550
rect -65 465 -55 535
rect -35 465 -20 535
rect -65 450 -20 465
rect -5 535 50 550
rect -5 465 10 535
rect 35 465 50 535
rect -5 450 50 465
rect 65 535 115 550
rect 65 465 80 535
rect 100 465 115 535
rect 65 450 115 465
rect 130 745 165 845
rect 180 830 230 845
rect 180 760 195 830
rect 215 760 230 830
rect 180 745 230 760
rect 130 550 155 745
rect 130 450 165 550
rect 180 535 230 550
rect 180 465 195 535
rect 215 465 230 535
rect 180 450 230 465
<< ndiffc >>
rect -55 300 -35 370
rect -55 0 -35 70
rect 65 300 85 370
rect 130 300 150 370
rect 195 300 215 370
rect 65 0 85 70
rect 130 0 150 70
rect 195 0 215 70
<< pdiffc >>
rect -55 760 -35 830
rect 10 760 35 830
rect 80 760 100 830
rect -55 465 -35 535
rect 10 465 35 535
rect 80 465 100 535
rect 195 760 215 830
rect 195 465 215 535
<< psubdiff >>
rect 130 -60 230 -45
rect 130 -80 145 -60
rect 215 -80 230 -60
rect 130 -95 230 -80
<< nsubdiff >>
rect 15 910 115 925
rect 15 890 30 910
rect 100 890 115 910
rect 15 875 115 890
<< psubdiffcont >>
rect 145 -80 215 -60
<< nsubdiffcont >>
rect 30 890 100 910
<< poly >>
rect -20 845 -5 860
rect 50 845 65 860
rect 115 845 130 860
rect 165 845 180 860
rect -20 550 -5 745
rect 50 710 65 745
rect 35 700 75 710
rect 35 680 45 700
rect 65 680 75 700
rect 35 670 75 680
rect 35 635 75 645
rect 35 615 45 635
rect 65 615 75 635
rect 35 605 75 615
rect 50 550 65 605
rect 165 730 180 745
rect 165 720 225 730
rect 165 715 195 720
rect 185 700 195 715
rect 215 700 225 720
rect 185 690 225 700
rect 165 655 210 665
rect 165 635 180 655
rect 200 635 210 655
rect 165 625 210 635
rect 165 550 180 625
rect -20 385 -5 450
rect 50 415 65 450
rect 115 415 130 450
rect 35 400 65 415
rect 100 400 130 415
rect 35 385 50 400
rect 100 385 115 400
rect 165 385 180 450
rect 35 245 50 285
rect 35 235 75 245
rect 35 215 45 235
rect 65 215 75 235
rect 35 205 75 215
rect 35 170 75 180
rect 35 150 45 170
rect 65 150 75 170
rect 35 140 75 150
rect 35 85 50 140
rect 100 85 115 285
rect 165 270 180 285
rect 165 260 220 270
rect 165 240 190 260
rect 210 240 220 260
rect 165 230 220 240
rect 140 180 180 190
rect 140 160 150 180
rect 170 160 180 180
rect 140 150 180 160
rect 165 85 180 150
rect -20 -55 -5 -15
rect 35 -30 50 -15
rect 100 -55 115 -15
rect 165 -30 180 -15
rect -20 -70 115 -55
rect -20 -115 20 -70
rect -20 -135 -10 -115
rect 10 -135 20 -115
rect -20 -145 20 -135
<< polycont >>
rect 45 680 65 700
rect 45 615 65 635
rect 195 700 215 720
rect 180 635 200 655
rect 45 215 65 235
rect 45 150 65 170
rect 190 240 210 260
rect 150 160 170 180
rect -10 -135 10 -115
<< locali >>
rect 20 910 110 920
rect 20 890 30 910
rect 100 890 110 910
rect 20 880 110 890
rect -85 830 -25 840
rect -85 760 -55 830
rect -35 760 -25 830
rect -85 750 -25 760
rect -5 830 45 840
rect -5 760 10 830
rect 35 760 45 830
rect -5 750 45 760
rect 70 830 110 880
rect 70 760 80 830
rect 100 760 110 830
rect 185 830 250 840
rect 185 770 195 830
rect 70 750 110 760
rect 145 760 195 770
rect 215 760 250 830
rect 145 750 250 760
rect -5 645 15 750
rect 35 700 75 710
rect 35 680 45 700
rect 65 690 75 700
rect 65 680 120 690
rect 35 670 120 680
rect -5 635 75 645
rect -5 625 45 635
rect 35 615 45 625
rect 65 615 75 635
rect 35 605 75 615
rect 100 585 120 670
rect 145 665 165 750
rect 185 720 225 730
rect 185 700 195 720
rect 215 710 225 720
rect 215 700 250 710
rect 185 690 250 700
rect 145 655 210 665
rect 145 635 180 655
rect 200 635 210 655
rect 145 625 210 635
rect 25 565 120 585
rect 25 545 45 565
rect 230 545 250 690
rect -85 535 -25 545
rect -85 465 -55 535
rect -35 465 -25 535
rect -85 455 -25 465
rect 0 535 45 545
rect 0 465 10 535
rect 35 465 45 535
rect 0 455 45 465
rect 70 535 110 545
rect 70 465 80 535
rect 100 465 110 535
rect 185 535 250 545
rect 185 475 195 535
rect 70 455 110 465
rect 140 465 195 475
rect 215 465 250 535
rect 140 455 250 465
rect 25 380 45 455
rect 140 380 160 455
rect -85 370 -25 380
rect -85 300 -55 370
rect -35 300 -25 370
rect 25 370 95 380
rect 25 360 65 370
rect 55 310 65 360
rect -85 290 -25 300
rect -5 300 65 310
rect 85 300 95 370
rect -5 290 95 300
rect 120 370 160 380
rect 120 300 130 370
rect 150 300 160 370
rect 120 290 160 300
rect 185 370 250 380
rect 185 300 195 370
rect 215 300 250 370
rect 185 290 250 300
rect -5 160 15 290
rect 35 235 75 245
rect 35 215 45 235
rect 65 225 75 235
rect 65 215 115 225
rect 35 205 115 215
rect 35 170 75 180
rect 35 160 45 170
rect -5 150 45 160
rect 65 150 75 170
rect -5 140 75 150
rect 95 120 115 205
rect 140 190 160 290
rect 180 260 220 270
rect 180 240 190 260
rect 210 240 220 260
rect 180 230 220 240
rect 140 180 180 190
rect 140 160 150 180
rect 170 160 180 180
rect 140 150 180 160
rect 200 130 220 230
rect 75 100 115 120
rect 140 110 220 130
rect 75 85 95 100
rect -85 70 -25 80
rect -85 0 -55 70
rect -35 0 -25 70
rect -85 -10 -25 0
rect 55 70 95 85
rect 140 80 160 110
rect 55 0 65 70
rect 85 0 95 70
rect 55 -10 95 0
rect 120 70 160 80
rect 120 0 130 70
rect 150 0 160 70
rect 120 -10 160 0
rect 185 70 250 80
rect 185 0 195 70
rect 215 0 250 70
rect 185 -10 250 0
rect 185 -50 225 -10
rect 135 -60 225 -50
rect 135 -80 145 -60
rect 215 -80 225 -60
rect 135 -90 225 -80
rect -20 -115 20 -105
rect -20 -135 -10 -115
rect 10 -135 20 -115
rect -20 -145 20 -135
<< viali >>
rect 30 890 100 910
rect 80 760 100 830
rect 80 465 100 535
rect -55 300 -35 370
rect 195 300 215 370
rect -55 0 -35 70
rect 195 0 215 70
rect 145 -80 215 -60
rect -10 -135 10 -115
<< metal1 >>
rect 20 910 110 920
rect 20 890 30 910
rect 100 890 110 910
rect 20 840 110 890
rect -85 830 250 840
rect -85 760 80 830
rect 100 760 250 830
rect -85 750 250 760
rect 70 535 110 750
rect 70 465 80 535
rect 100 465 110 535
rect 70 455 110 465
rect -85 370 -25 380
rect -85 300 -55 370
rect -35 300 -25 370
rect -85 290 -25 300
rect -65 80 -25 290
rect 185 370 250 380
rect 185 300 195 370
rect 215 300 250 370
rect 185 290 250 300
rect 185 80 225 290
rect -85 70 250 80
rect -85 0 -55 70
rect -35 0 195 70
rect 215 0 250 70
rect -85 -10 250 0
rect 135 -60 225 -10
rect 135 -80 145 -60
rect 215 -80 225 -60
rect 135 -90 225 -80
rect -85 -115 250 -105
rect -85 -135 -10 -115
rect 10 -135 250 -115
rect -85 -145 250 -135
<< labels >>
rlabel locali -85 795 -85 795 7 D
port 2 w
rlabel locali -85 500 -85 500 7 Dn
port 4 w
rlabel locali 250 500 250 500 3 Qn
port 5 e
rlabel locali 250 795 250 795 3 Q
port 3 e
rlabel metal1 -85 35 -85 35 7 VN
port 6 w
rlabel metal1 -85 -125 -85 -125 7 CLK
port 7 w
rlabel metal1 -85 795 -85 795 7 VP
port 1 w
<< end >>
