magic
tech sky130A
timestamp 1695876091
<< error_p >>
rect 25 100 90 125
rect 0 0 50 100
rect 65 0 115 100
rect 25 -25 90 0
<< nmos >>
rect 50 0 65 100
<< ndiff >>
rect 0 0 50 100
rect 65 0 115 100
<< end >>
